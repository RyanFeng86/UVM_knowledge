`include "uvm_macros.svh"  
`include "transaction_write.sv"
import uvm_pkg::*; 

typedef uvm_sequencer #(my_write_transaction) my_write_sequencer;

