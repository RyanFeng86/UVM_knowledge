`ifndef sequencer_write_SV
`define sequencer_write_SV

`include "transaction_write.sv"


typedef uvm_sequencer #(my_write_transaction) my_write_sequencer;
`endif
