`ifndef testcase_da3_SV
`define testcase_da3_SV

`include "env.sv"
`include "sequence.sv"
`include "transaction_da3.sv"
`include "testcase.sv"

class my_test_da3 extends my_test;
    `uvm_component_utils(my_test_da3)

    function new(string name="",uvm_component parent);
        super.new(name,parent);
    endfunction

    virtual function void build_phase(uvm_phase phase);
        super.build_phase(phase);
        set_type_override_by_type(my_transaction::get_type(),my_transaction_da3::get_type()); //use factory replace/override my_transaction with my_transaction_da3
    endfunction

    virtual function void report_phase(uvm_phase phase);
        super.report_phase(phase);
        factory.print();//printed information in the log file start from factory configuration block. It shows orignal override to which targeting type
    endfunction

endclass



`endif