`ifndef sequencer_read_SV
`define sequencer_read_SV
 
`include "transaction_read.sv"


typedef uvm_sequencer #(my_read_transaction) my_read_sequencer;
`endif
