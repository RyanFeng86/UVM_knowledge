program automatic test;
    `include "testcase.sv"

    initial begin
        run_test();
    end
endprogram
